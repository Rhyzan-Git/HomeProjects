--Notes:
